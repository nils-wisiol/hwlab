`timescale 1ns / 1ps
module PinGen(
    input wire clk,
    input wire en,
    output reg [] counter,
    output reg [] pin
    );


endmodule
