`timescale 1ns / 1ps

module Ex11_tb();

reg tb_a;
reg tb_b;
wire tb_s;
wire tb_c;

Ex11 andi(
	.A(tb_a),
	.B(tb_b),
	.S(tb_s),
	.C(tb_c));

initial
begin
	tb_a <= 1'b0;  // 1 bit, value zero
	tb_b <= 1'b0;
end

always
begin
	#50 tb_a <= ~tb_a;
end

always
begin
	#100 tb_b <= ~tb_b;
end

endmodule
